
// Global Params 
`define NUM_STAGES 15
`define KDCO_COARSE 250e6
`define KDCO_FINE 10e5 

