
// Global Params 
`define NUM_STAGES 15
`define REFCLK_PERIOD 8*1000*1000
`define KDCO_COARSE 250e6
`define KDCO_FINE 1e4 //50e6

