`timescale 1fs/1fs


module dco (
    input  int dctrl_coarse,
    input  int dctrl_fine,
    input  logic refclk,
    input  logic resetn,
    output logic pclk, 
    output int dco_phase
);
    // DCO I/O Interface

endmodule

