`timescale 1fs/1fs


module pd (
    input  logic refclk,
    input  logic fbclk,
    input  logic resetn,
    output int out
);
    // hase Detector IO

endmodule

